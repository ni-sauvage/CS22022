----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 28.12.2021 01:05:12
-- Design Name: 
-- Module Name: Control_Memory42Bit_256_20334203 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Control_Memory42Bit_256_InitTB_20334203 is
    Port (IN_CAR : in std_logic_vector(16 downto 0);
        FL : out std_logic; -- 0
        RZ : out std_logic; -- 1
        RN : out std_logic; -- 2
        RC : out std_logic; -- 3
        RV : out std_logic; -- 4
        MW : out std_logic; -- 5
        MM : out std_logic; -- 6
        RW : out std_logic; -- 7
        MD : out std_logic; -- 8
        FS : out std_logic_vector(4 downto 0); -- 9 to 13
        MB : out std_logic; -- 14
        TB : out std_logic; -- 15
        TA : out std_logic; -- 16
        TD : out std_logic; -- 17
        PL : out std_logic; -- 18
        PI : out std_logic; -- 19
        IL : out std_logic; -- 20
        MC : out std_logic; -- 21
        MS : out std_logic_vector(2 downto 0); -- 22 to 24
        NA : out std_logic_vector(16 downto 0) -- 25 to 41
    );
end Control_Memory42Bit_256_InitTB_20334203;

architecture Behavioral of Control_Memory42Bit_256_InitTB_20334203 is

type mem_array is array(0 to 255) of std_logic_vector(41 downto 0);
-- initialise the control memory
signal control_mem : mem_array := (
-- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
-- | Next Address | MS | M| I| P| P| T| T| T| M| FS |M|R|M|M|R|R|R|R|F|
-- | Next Address | MS | C| L| I| L| D| A| B| B| FS |D|W|M|W|V|C|N|Z|L|
-- "00000000000000000 000 0 0 0 0 0 0 0 0 00000 0 0 0 0 0 0 0 0 0"
    "000000000000000000000000000000000000000011",
    "000000000000000000000000000000000000000100",
    "000000000000000000000000000000000000000101",
    "000000000000000000000000000000000000000110",
    "000000000000000000000000000000000000000111",
    "000000000000000000000000000000000000001000",
    "000000000000000000000000000000000000001001",
    "000000000000000000000000000000000000001010",
    "000000000000000000000000000000000000001011",
    "000000000000000000000000000000000000001100",
    "000000000000000000000000000000000000001101",
    "000000000000000000000000000000000000001110",
    "000000000000000000000000000000000000001111",
    "000000000000000000000000000000000000010000",
    "000000000000000000000000000000000000010001",
    "000000000000000000000000000000000000010010",
    "000000000000000000000000000000000000010011",
    "000000000000000000000000000000000000010100",
    "000000000000000000000000000000000000010101",
    "000000000000000000000000000000000000010110",
    "000000000000000000000000000000000000010111",
    "000000000000000000000000000000000000011000",
    "000000000000000000000000000000000000011001",
    "000000000000000000000000000000000000011010",
    "000000000000000000000000000000000000011011",
    "000000000000000000000000000000000000011100",
    "000000000000000000000000000000000000011101",
    "000000000000000000000000000000000000011110",
    "000000000000000000000000000000000000011111",
    "000000000000000000000000000000000000100000",
    "000000000000000000000000000000000000100001",
    "000000000000000000000000000000000000100010",
    "000000000000000000000000000000000000100011",
    "000000000000000000000000000000000000100100",
    "000000000000000000000000000000000000100101",
    "000000000000000000000000000000000000100110",
    "000000000000000000000000000000000000100111",
    "000000000000000000000000000000000000101000",
    "000000000000000000000000000000000000101001",
    "000000000000000000000000000000000000101010",
    "000000000000000000000000000000000000101011",
    "000000000000000000000000000000000000101100",
    "000000000000000000000000000000000000101101",
    "000000000000000000000000000000000000101110",
    "000000000000000000000000000000000000101111",
    "000000000000000000000000000000000000110000",
    "000000000000000000000000000000000000110001",
    "000000000000000000000000000000000000110010",
    "000000000000000000000000000000000000110011",
    "000000000000000000000000000000000000110100",
    "000000000000000000000000000000000000110101",
    "000000000000000000000000000000000000110110",
    "000000000000000000000000000000000000110111",
    "000000000000000000000000000000000000111000",
    "000000000000000000000000000000000000111001",
    "000000000000000000000000000000000000111010",
    "000000000000000000000000000000000000111011",
    "000000000000000000000000000000000000111100",
    "000000000000000000000000000000000000111101",
    "000000000000000000000000000000000000111110",
    "000000000000000000000000000000000000111111",
    "000000000000000000000000000000000001000000",
    "000000000000000000000000000000000001000001",
    "000000000000000000000000000000000001000010",
    "000000000000000000000000000000000001000011",
    "000000000000000000000000000000000001000100",
    "000000000000000000000000000000000001000101",
    "000000000000000000000000000000000001000110",
    "000000000000000000000000000000000001000111",
    "000000000000000000000000000000000001001000",
    "000000000000000000000000000000000001001001",
    "000000000000000000000000000000000001001010",
    "000000000000000000000000000000000001001011",
    "000000000000000000000000000000000001001100",
    "000000000000000000000000000000000001001101",
    "000000000000000000000000000000000001001110",
    "000000000000000000000000000000000001001111",
    "000000000000000000000000000000000001010000",
    "000000000000000000000000000000000001010001",
    "000000000000000000000000000000000001010010",
    "000000000000000000000000000000000001010011",
    "000000000000000000000000000000000001010100",
    "000000000000000000000000000000000001010101",
    "000000000000000000000000000000000001010110",
    "000000000000000000000000000000000001010111",
    "000000000000000000000000000000000001011000",
    "000000000000000000000000000000000001011001",
    "000000000000000000000000000000000001011010",
    "000000000000000000000000000000000001011011",
    "000000000000000000000000000000000001011100",
    "000000000000000000000000000000000001011101",
    "000000000000000000000000000000000001011110",
    "000000000000000000000000000000000001011111",
    "000000000000000000000000000000000001100000",
    "000000000000000000000000000000000001100001",
    "000000000000000000000000000000000001100010",
    "000000000000000000000000000000000001100011",
    "000000000000000000000000000000000001100100",
    "000000000000000000000000000000000001100101",
    "000000000000000000000000000000000001100110",
    "000000000000000000000000000000000001100111",
    "000000000000000000000000000000000001101000",
    "000000000000000000000000000000000001101001",
    "000000000000000000000000000000000001101010",
    "000000000000000000000000000000000001101011",
    "000000000000000000000000000000000001101100",
    "000000000000000000000000000000000001101101",
    "000000000000000000000000000000000001101110",
    "000000000000000000000000000000000001101111",
    "000000000000000000000000000000000001110000",
    "000000000000000000000000000000000001110001",
    "000000000000000000000000000000000001110010",
    "000000000000000000000000000000000001110011",
    "000000000000000000000000000000000001110100",
    "000000000000000000000000000000000001110101",
    "000000000000000000000000000000000001110110",
    "000000000000000000000000000000000001110111",
    "000000000000000000000000000000000001111000",
    "000000000000000000000000000000000001111001",
    "000000000000000000000000000000000001111010",
    "000000000000000000000000000000000001111011",
    "000000000000000000000000000000000001111100",
    "000000000000000000000000000000000001111101",
    "000000000000000000000000000000000001111110",
    "000000000000000000000000000000000001111111",
    "000000000000000000000000000000000010000000",
    "000000000000000000000000000000000010000001",
    "000000000000000000000000000000000010000010",
    "000000000000000000000000000000000010000011",
    "000000000000000000000000000000000010000100",
    "000000000000000000000000000000000010000101",
    "000000000000000000000000000000000010000110",
    "000000000000000000000000000000000010000111",
    "000000000000000000000000000000000010001000",
    "000000000000000000000000000000000010001001",
    "000000000000000000000000000000000010001010",
    "000000000000000000000000000000000010001011",
    "000000000000000000000000000000000010001100",
    "000000000000000000000000000000000010001101",
    "000000000000000000000000000000000010001110",
    "000000000000000000000000000000000010001111",
    "000000000000000000000000000000000010010000",
    "000000000000000000000000000000000010010001",
    "000000000000000000000000000000000010010010",
    "000000000000000000000000000000000010010011",
    "000000000000000000000000000000000010010100",
    "000000000000000000000000000000000010010101",
    "000000000000000000000000000000000010010110",
    "000000000000000000000000000000000010010111",
    "000000000000000000000000000000000010011000",
    "000000000000000000000000000000000010011001",
    "000000000000000000000000000000000010011010",
    "000000000000000000000000000000000010011011",
    "000000000000000000000000000000000010011100",
    "000000000000000000000000000000000010011101",
    "000000000000000000000000000000000010011110",
    "000000000000000000000000000000000010011111",
    "000000000000000000000000000000000010100000",
    "000000000000000000000000000000000010100001",
    "000000000000000000000000000000000010100010",
    "000000000000000000000000000000000010100011",
    "000000000000000000000000000000000010100100",
    "000000000000000000000000000000000010100101",
    "000000000000000000000000000000000010100110",
    "000000000000000000000000000000000010100111",
    "000000000000000000000000000000000010101000",
    "000000000000000000000000000000000010101001",
    "000000000000000000000000000000000010101010",
    "000000000000000000000000000000000010101011",
    "000000000000000000000000000000000010101100",
    "000000000000000000000000000000000010101101",
    "000000000000000000000000000000000010101110",
    "000000000000000000000000000000000010101111",
    "000000000000000000000000000000000010110000",
    "000000000000000000000000000000000010110001",
    "000000000000000000000000000000000010110010",
    "000000000000000000000000000000000010110011",
    "000000000000000000000000000000000010110100",
    "000000000000000000000000000000000010110101",
    "000000000000000000000000000000000010110110",
    "000000000000000000000000000000000010110111",
    "000000000000000000000000000000000010111000",
    "000000000000000000000000000000000010111001",
    "000000000000000000000000000000000010111010",
    "000000000000000000000000000000000010111011",
    "000000000000000000000000000000000010111100",
    "000000000000000000000000000000000010111101",
    "000000000000000000000000000000000010111110",
    "000000000000000000000000000000000010111111",
    "000000000000000000000000000000000011000000",
    "000000000000000000000000000000000011000001",
    "000000000000000000000000000000000011000010",
    "000000000000000000000000000000000011000011",
    "000000000000000000000000000000000011000100",
    "000000000000000000000000000000000011000101",
    "000000000000000000000000000000000011000110",
    "000000000000000000000000000000000011000111",
    "000000000000000000000000000000000011001000",
    "000000000000000000000000000000000011001001",
    "000000000000000000000000000000000011001010",
    "000000000000000000000000000000000011001011",
    "000000000000000000000000000000000011001100",
    "000000000000000000000000000000000011001101",
    "000000000000000000000000000000000011001110",
    "000000000000000000000000000000000011001111",
    "000000000000000000000000000000000011010000",
    "000000000000000000000000000000000011010001",
    "000000000000000000000000000000000011010010",
    "000000000000000000000000000000000011010011",
    "000000000000000000000000000000000011010100",
    "000000000000000000000000000000000011010101",
    "000000000000000000000000000000000011010110",
    "000000000000000000000000000000000011010111",
    "000000000000000000000000000000000011011000",
    "000000000000000000000000000000000011011001",
    "000000000000000000000000000000000011011010",
    "000000000000000000000000000000000011011011",
    "000000000000000000000000000000000011011100",
    "000000000000000000000000000000000011011101",
    "000000000000000000000000000000000011011110",
    "000000000000000000000000000000000011011111",
    "000000000000000000000000000000000011100000",
    "000000000000000000000000000000000011100001",
    "000000000000000000000000000000000011100010",
    "000000000000000000000000000000000011100011",
    "000000000000000000000000000000000011100100",
    "000000000000000000000000000000000011100101",
    "000000000000000000000000000000000011100110",
    "000000000000000000000000000000000011100111",
    "000000000000000000000000000000000011101000",
    "000000000000000000000000000000000011101001",
    "000000000000000000000000000000000011101010",
    "000000000000000000000000000000000011101011",
    "000000000000000000000000000000000011101100",
    "000000000000000000000000000000000011101101",
    "000000000000000000000000000000000011101110",
    "000000000000000000000000000000000011101111",
    "000000000000000000000000000000000011110000",
    "000000000000000000000000000000000011110001",
    "000000000000000000000000000000000011110010",
    "000000000000000000000000000000000011110011",
    "000000000000000000000000000000000011110100",
    "000000000000000000000000000000000011110101",
    "000000000000000000000000000000000011110110",
    "000000000000000000000000000000000011110111",
    "000000000000000000000000000000000011111000",
    "000000000000000000000000000000000011111001",
    "000000000000000000000000000000000011111010",
    "000000000000000000000000000000000011111011",
    "000000000000000000000000000000000011111100",
    "000000000000000000000000000000000011111101",
    "000000000000000000000000000000000011111110",
    "000000000000000000000000000000000011111111",
    "000000000000000000000000000000000100000000",
    "000000000000000000000000000000000100000001",
    "000000000000000000000000000000000100000010"

    );                                                          
signal content_at_address : std_logic_vector(41 downto 0);
begin
    content_at_address <= control_mem(to_integer(unsigned(IN_CAR(8 downto 0)))) after 2ns;
    FL <= content_at_address(0); -- 0
    RZ <= content_at_address(1); -- 1
    RN <= content_at_address(2); -- 2
    RC <= content_at_address(3); -- 3
    RV <= content_at_address(4); -- 4
    MW <= content_at_address(5); -- 5
    MM <= content_at_address(6); -- 6
    RW <= content_at_address(7); -- 7
    MD <= content_at_address(8); -- 8
    FS <= content_at_address(13 downto 9); -- 9 to 13
    MB <= content_at_address(14); -- 14
    TB <= content_at_address(15); -- 15
    TA <= content_at_address(16); -- 16
    TD <= content_at_address(17); -- 17
    PL <= content_at_address(18); -- 18
    PI <= content_at_address(19); -- 19
    IL <= content_at_address(20); -- 20
    MC <= content_at_address(21); -- 21
    MS <= content_at_address(24 downto 22); -- 22 to 24
    NA <= content_at_address(41 downto 25); -- 25 to 41

end Behavioral;
